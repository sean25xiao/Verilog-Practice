module top_module ( input a, input b, output out );

    mod_a my_module ( .in1(a), .in2(b), .out(out), );

endmodule
